module basic(out, a, b);

output [2:0] out;
input [2:0] a;
input [2:0] b;

assign out = a + b;

endmodule
