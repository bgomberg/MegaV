`ifndef __MEM_OP_SIZE_SV__
`define __MEM_OP_SIZE_SV__

`define MEM_OP_SIZE_BYTE 2'b00
`define MEM_OP_SIZE_HALF_WORD 2'b01
`define MEM_OP_SIZE_WORD 2'b10

`endif
