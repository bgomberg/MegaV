`ifndef __FSM_FAULT_NUM_SV__
`define __FSM_FAULT_NUM_SV__

`define FSM_FAULT_NUM_INSTR_ADDR_MISALIGNED 3'b000
`define FSM_FAULT_NUM_INSTR_ACCESS_FAULT 3'b001
`define FSM_FAULT_NUM_ILLEGAL_INSTR 3'b010
`define FSM_FAULT_NUM_LOAD_ADDR_MISALIGNED 3'b100
`define FSM_FAULT_NUM_LOAD_ACCESS_FAULT 3'b101
`define FSM_FAULT_NUM_STORE_ADDR_MISALIGNED 3'b110
`define FSM_FAULT_NUM_STORE_ACCESS_FAULT 3'b111

`endif
