`ifndef __FSM_FAULT_NUM_SV__
`define __FSM_FAULT_NUM_SV__

`define MEM_FAULT_NUM_LOAD_ADDR_MISALIGNED 2'b00
`define MEM_FAULT_NUM_LOAD_ACCESS_FAULT 2'b01
`define MEM_FAULT_NUM_STORE_ADDR_MISALIGNED 2'b10
`define MEM_FAULT_NUM_STORE_ACCESS_FAULT 2'b11

`endif
