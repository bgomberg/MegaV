`include "cells/dff.sv"
`include "cells/dff_stages.sv"
`include "cells/dffe.sv"
`include "cells/mux2.sv"
`include "cells/mux4.sv"
`include "constants/fsm_control_op.sv"
`include "constants/fsm_fault_num.sv"
`include "constants/stages.sv"

/*
 * FSM.
 */
module fsm(
    input logic clk, // Clock signal
    input logic reset_n, // Reset signal (active low)
    input logic illegal_instr_fault, // Illegal instruction fault
    input logic [2:0] mem_fault_num, // Memory fault number
    input logic ext_int, // External interrupt
    input logic sw_int, // Software interrupt
    output logic [`NUM_STAGES-1:0] stage_active_n, // Current stage (active low)
    output logic [1:0] control_op, // Control operation
    output logic [2:0] fault_num // Active fault number
);

    /* Next Stage */
    wire [`NUM_STAGES-1:0] next_stage_n = {stage_active_n[`NUM_STAGES-2:0], stage_active_n[`NUM_STAGES-1]};

    /* In Progress */
    logic in_progress;
    dff in_progress_dff(
        .clk(clk),
        .clear_n(reset_n),
        .in(~in_progress),
        .out(in_progress)
    );

    /* Control Op */
    wire fault_value;
    mux2 fault_value_mux(
        .a(fault),
        .b(active_fault),
        .select(in_progress),
        .out(fault_value)
    );
    wire [1:0] control_op_value = {~fault_value & ~ext_int, ~fault_value & (ext_int | ~sw_int)};
    // TODO: There are some weird bugs that get exposed if this signal is simplified or non-public
    wire update_control_op /* verilator public */ = ~reset_n | (in_progress & (~next_stage_n[`STAGE_CONTROL] | active_fault));
    dffe #(.BITS(2)) control_op_dffe(
        .clk(clk),
        .clear_n(reset_n),
        .enable_n(~update_control_op),
        .in(control_op_value),
        .out(control_op)
    );

    /* Fault / Fault Number */
    logic fault;
    wire mem_fault = mem_fault_num[2];
    wire fetch_stage_mem_fault = mem_fault & ~stage_active_n[`STAGE_FETCH];
    wire mem_stage_mem_fault = mem_fault & ~stage_active_n[`STAGE_MEMORY];
    wire non_control_stage_instr_fault = stage_active_n[`STAGE_CONTROL] & illegal_instr_fault;
    wire active_fault = in_progress & (fetch_stage_mem_fault | mem_stage_mem_fault | non_control_stage_instr_fault);
    wire [2:0] next_fault_num = {
        mem_stage_mem_fault & ~non_control_stage_instr_fault,
        (mem_stage_mem_fault & mem_fault_num[1]) | non_control_stage_instr_fault,
        ~non_control_stage_instr_fault & mem_fault_num[0]
    };
    dffe fault_dff(
        .clk(clk),
        .clear_n(reset_n),
        .enable_n(~in_progress),
        .in(active_fault),
        .out(fault)
    );
    dffe #(.BITS(3)) fault_num_dffe(
        .clk(clk),
        .clear_n(reset_n),
        .enable_n(~active_fault),
        .in(next_fault_num),
        .out(fault_num)
    );

    /* Active Stage */
    wire [`NUM_STAGES-1:0] next_stage_active_n;
    mux4 #(.BITS(`NUM_STAGES)) next_stage_active_n_mux(
        .d1(stage_active_n),
        .d2(stage_active_n),
        .d3(next_stage_n),
        .d4(~`DEFAULT_STAGE_ACTIVE),
        .select({in_progress, active_fault}),
        .out(next_stage_active_n)
    );
    dff_stages stage_active_dff(
        .clk(clk),
        .clear_n(reset_n),
        .in(next_stage_active_n),
        .out(stage_active_n)
    );

`ifdef FORMAL
    initial assume(~reset_n);
    logic f_past_valid;
    initial f_past_valid = 0;
    always_ff @(posedge clk) begin
        f_past_valid = 1;
    end

    /* Validate logic */
    wire [`NUM_STAGES-1:0] stage_active = ~stage_active_n;
    always_ff @(posedge clk) begin
        if (f_past_valid) begin
            // Only one bit in stage_active should ever be set
            assume($past(stage_active & (stage_active - 1)) == 0);
            if ($past(~reset_n)) begin
                assert(stage_active == 1 << 0);
            end else if ($past(stage_active) != $past(stage_active, 2) || $past(~reset_n, 2)) begin
                // need to stay in each stage for at least 2 clock cycles
                assert(stage_active == $past(stage_active));
            end else begin
                assert(stage_active == (1 << 0) || stage_active != $past(stage_active));
                if ($past(illegal_instr_fault) && !$past(stage_active[`STAGE_CONTROL])) begin
                    assert(stage_active == (1 << 0));
                    assert(fault_num == `FSM_FAULT_NUM_ILLEGAL_INSTR);
                end else if ($past(mem_fault_num[2] & ~mem_fault_num[0]) && $past(stage_active[`STAGE_FETCH])) begin
                    assert(stage_active == (1 << 0));
                    assert(fault_num == `FSM_FAULT_NUM_INSTR_ADDR_MISALIGNED);
                end else if ($past(mem_fault_num[2] & ~mem_fault_num[0]) && $past(stage_active[`STAGE_MEMORY])) begin
                    assert(stage_active == (1 << 0));
                    if ($past(mem_fault_num[1])) begin
                        assert(fault_num == `FSM_FAULT_NUM_STORE_ADDR_MISALIGNED);
                    end else begin
                        assert(fault_num == `FSM_FAULT_NUM_LOAD_ADDR_MISALIGNED);
                    end
                end else if ($past(mem_fault_num[2] & mem_fault_num[0]) && $past(stage_active[`STAGE_FETCH])) begin
                    assert(fault_num == `FSM_FAULT_NUM_INSTR_ACCESS_FAULT);
                end else if ($past(mem_fault_num[2] & mem_fault_num[0]) && $past(stage_active[`STAGE_MEMORY])) begin
                    assert(stage_active == (1 << 0));
                    if ($past(mem_fault_num[1])) begin
                        assert(fault_num == `FSM_FAULT_NUM_STORE_ACCESS_FAULT);
                    end else begin
                        assert(fault_num == `FSM_FAULT_NUM_LOAD_ACCESS_FAULT);
                    end
                end else begin
                    // Stage was completed without a fault
                    assert(stage_active == $past({stage_active[`NUM_STAGES-2:0], stage_active[`NUM_STAGES-1]}));
                end
            end
        end
    end
`endif

endmodule
