`ifndef __ALU_MICROCODE_SV__
`define __ALU_MICROCODE_SV__

`include "types.sv"

`define ALU_MICROCODE_ADD               {4'b0000, SHIFTER_OP_SLL, ALU_OUTPUT_SELECT_ADD_SUB}
`define ALU_MICROCODE_SUB               {4'b0001, SHIFTER_OP_SLL, ALU_OUTPUT_SELECT_ADD_SUB}
`define ALU_MICROCODE_SLL               {4'b0000, SHIFTER_OP_SLL, ALU_OUTPUT_SELECT_SLL}
`define ALU_MICROCODE_SRL               {4'b0000, SHIFTER_OP_SRL, ALU_OUTPUT_SELECT_SRL_SRA}
`define ALU_MICROCODE_SRA               {4'b0000, SHIFTER_OP_SRA, ALU_OUTPUT_SELECT_SRL_SRA}
`define ALU_MICROCODE_SLT               {4'b0001, SHIFTER_OP_SLL, ALU_OUTPUT_SELECT_SLT_BRANCH}
`define ALU_MICROCODE_SLTU              {4'b0011, SHIFTER_OP_SLL, ALU_OUTPUT_SELECT_SLTU}
`define ALU_MICROCODE_BEQ               {4'b1001, SHIFTER_OP_SLL, ALU_OUTPUT_SELECT_SLT_BRANCH}
`define ALU_MICROCODE_BNE               {4'b1101, SHIFTER_OP_SLL, ALU_OUTPUT_SELECT_SLT_BRANCH}
`define ALU_MICROCODE_BLT               {4'b0001, SHIFTER_OP_SLL, ALU_OUTPUT_SELECT_SLT_BRANCH}
`define ALU_MICROCODE_BGE               {4'b0101, SHIFTER_OP_SLL, ALU_OUTPUT_SELECT_SLT_BRANCH}
`define ALU_MICROCODE_BLTU              {4'b0011, SHIFTER_OP_SLL, ALU_OUTPUT_SELECT_SLT_BRANCH}
`define ALU_MICROCODE_BGEU              {4'b0111, SHIFTER_OP_SLL, ALU_OUTPUT_SELECT_SLT_BRANCH}
`define ALU_MICROCODE_XOR               {4'b0000, SHIFTER_OP_SLL, ALU_OUTPUT_SELECT_XOR}
`define ALU_MICROCODE_OR                {4'b0000, SHIFTER_OP_SLL, ALU_OUTPUT_SELECT_OR}
`define ALU_MICROCODE_AND               {4'b0000, SHIFTER_OP_SLL, ALU_OUTPUT_SELECT_AND}

`endif
