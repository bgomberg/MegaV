`ifndef __CSR_OP_SV__
`define __CSR_OP_SV__

`define CSR_OP_EXCEPTION    3'b000
`define CSR_OP_MRET         3'b001
`define CSR_OP_NO_OP        3'b011
`define CSR_OP_CSRRW        3'b101
`define CSR_OP_CSRRS        3'b110
`define CSR_OP_CSRRC        3'b111

`endif
